module ROM(input clock, input [31:0] address, output reg [32:0] instruction);

    reg [31:0] rom [1023:0]; 
    integer i;
    initial begin 
	 	rom[0] = 32'b10000000000000010000011000001010;
	 	rom[1] = 32'b00000100000000010001000000000000;
	 	rom[2] = 32'b00001100000000010001100000000000;
	 	rom[3] = 32'b00010100010000110010000000000000;
	 	rom[4] = 32'b10000100011001010001101000110100;
	 	rom[5] = 32'b00011000011001000010100000000000;
	 	rom[6] = 32'b00011100101000000011000000000000;
	 	rom[7] = 32'b00011100100000000101100000000000;
	 	rom[8] = 32'b00001100101001010010100000000000;
	 	rom[9] = 32'b10000000000000010000010000000000;
	 	rom[10] = 32'b10010100001000100000000000000000;
	 	rom[11] =  32'b10010000001001010000000000000000;
    end 

    always @ (posedge clock)
    begin 
        instruction = rom[address];
    end 

endmodule 