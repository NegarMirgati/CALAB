module ID (
	input clock, 
	input reset, 
	input [31:0] instruction
);

	

endmodule