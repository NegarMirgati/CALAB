module ConditionCheck(
	input [31:0] val1, 
	input [31:0] src2_val, 
	input [1:0] branch_type, 
	output [31:0] branch_tacken
	);

endmodule