module ROM(input clock, input [31:0] address, output reg [32:0] instruction);

    reg [31:0] rom [1023:0]; 
    integer i;
    initial begin 
	 rom[0] = 32'b10000000000000010000011000001010;
	 rom[1] = 32'b000001_00000_00001_00010_00000000000;
	 rom[2] = 32'b000011_00000_00001_00011_00000000000;
	 rom[3] = 32'b000101_00010_00011_00100_00000000000;
	 rom[4] = 32'b100001_00011_00101_00011_01000110100;
	 rom[5] = 32'b000110_00011_00100_00101_00000000000;
	 rom[6] = 32'b000111_00101_00000_00110_00000000000;
	 rom[7] = 32'b000111_00100_00000_01011_00000000000;
	 rom[8] = 32'b000011_00101_00101_00101_00000000000;
	 rom[9] = 32'b100000_00000_00001_00000_10000000000;
	 rom[10] = 32'b100101_00001_00010_00000_00000000000;
	 rom[11] =  32'b100100_00001_00101_00000_00000000000;
	
    end 

    always @ (posedge clock)
    begin 
        instruction = rom[address];
    end 

endmodule 