module AddressMapping(
	input [31:0] input_val, 
	output [31:0] address
);
	
	// change later 
	assign address = input_val;

endmodule 