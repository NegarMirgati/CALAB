module MUX  #(parameter LEN = 32) (
);


endmodule 