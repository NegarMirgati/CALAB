module ROM(input clock,input reset, input [31:0] address, output [31:0] instruction);

    reg [7:0] rom [400:0]; 
    integer i;

    always @ (posedge clock) begin 
    if(reset) begin 
	  /*1*/	{rom[0], rom[1], rom[2], rom[3]} = 32'b10000000000000010000011000001010;
	 
	       	{rom[4], rom[5], rom[6], rom[7]} = 32'd0;
	        {rom[8], rom[9], rom[10], rom[11]} = 32'd0;
	 	
	 /*2*/ 	{rom[12], rom[13], rom[14], rom[15]} = 32'b00000100000000010001000000000000;

	 	
	 /*3*/ 	{rom[16], rom[17], rom[18], rom[19]} = 32'b00001100000000010001100000000000;
	 	
	       	{rom[20], rom[21], rom[22], rom[23]} = 32'd0;
	 	      {rom[24], rom[25], rom[26], rom[27]} = 32'd0;
	 	
	 /*4*/	{rom[28], rom[29], rom[30], rom[31]} = 32'b00010100010000110010000000000000;
	 /*5*/	{rom[32], rom[33], rom[34], rom[35]} = 32'b10000100011001010001101000110100;

	 /*6*/	{rom[36], rom[37], rom[38], rom[39]} = 32'b00011000011001000010100000000000;
	 
	 	 	
	   	   {rom[40], rom[41], rom[42], rom[43]} = 32'd0;
	 	     {rom[44], rom[45], rom[46], rom[47]} = 32'd0;
	 
	 	/* 7 */ {rom[48], rom[49], rom[50], rom[51]} = 32'b00011100101000000011000000000000;
	 	
	 	/* 8 */ {rom[52], rom[53], rom[54], rom[55]} = 32'b00011100100000000101100000000000;
	 	/* 9 */ {rom[56], rom[57], rom[58], rom[59]} = 32'b00001100101001010010100000000000;
	 	/* 10 */ {rom[60], rom[61], rom[62], rom[63]} = 32'b10000000000000010000010000000000;
	 	
	 	{rom[64], rom[65], rom[66], rom[67]} = 32'd0;
	 	{rom[68], rom[69], rom[70], rom[71]} = 32'd0;
	 	
	 	/* 11 */ {rom[72], rom[73], rom[74], rom[75]} = 32'b10010100001000100000000000000000;
	 	
	 	/* 12 */ {rom[76], rom[77], rom[78], rom[79]} =  32'b10010000001001010000000000000000;
	  
	  {rom[80], rom[81], rom[82], rom[83]} = 32'd0;
	 	{rom[84], rom[85], rom[86], rom[87]} = 32'd0;
	 	
	 
    /* 13 */ {rom[88], rom[89], rom[90], rom[91]} = 32'b10100000101000000000000000000001; 
     /* 14 */ {rom[92], rom[93], rom[94], rom[95]}  = 32'b00100000101000010011100000000000;
     /* 15 */{ rom[96], rom[97], rom[98], rom[99]} =  32'b001000_00101_00001_00000_00000000000;
    /* 16 */ { rom[100], rom[101], rom[102], rom[103]} = 32'b001001_00011_01011_00111_00000000000;
    /* 17 */ { rom[104], rom[105], rom[106], rom[107]} = 32'b001010_00011_01011_01000_00000000000;
    /* 18 */ { rom[108], rom[109], rom[110], rom[111]} = 32'b001011_00011_00100_01001_00000000000;
    /* 19 */ { rom[112], rom[113], rom[114], rom[115]} = 32'b001100_00011_00100_01010_00000000000;
    /* 20 */ { rom[116], rom[117], rom[118], rom[119]} = 32'b100101_00001_00011_00000_00000000100;
    /* 21 */ { rom[120], rom[121], rom[122], rom[123]} = 32'b100101_00001_00100_00000_00000001000;
    /* 22 */ { rom[124], rom[125], rom[126], rom[127]} = 32'b100101_00001_00101_00000_00000001100;
    /* 23 */ { rom[128], rom[129], rom[130], rom[131]} = 32'b100101_00001_00110_00000_00000010000;
    /* 24 */ { rom[132], rom[133], rom[134], rom[135]} = 32'b100100_00001_01011_00000_00000000100;
    /* 25 */ { rom[136], rom[137], rom[138], rom[139]} =32'b100101_00001_00111_00000_00000010100; 
    /* 26 */ { rom[140], rom[141], rom[142], rom[143]} = 32'b100101_00001_01000_00000_00000011000;
    /* 27 */ { rom[144], rom[145], rom[146], rom[147]} = 32'b100101_00001_01001_00000_00000011100;
    /* 28 */ { rom[148], rom[149], rom[150], rom[151]} = 32'b100101_00001_01010_00000_00000100000;
    /* 29 */ { rom[152], rom[153], rom[154], rom[155]} = 32'b100101_00001_01011_00000_00000100100;
    /* 30 */ { rom[156], rom[157], rom[158], rom[159]} = 32'b100000_00000_00001_00000_00000000011;
    /* 31 */ { rom[160], rom[161], rom[162], rom[163]} = 32'b100000_00000_00100_00000_10000000000;


  /* 32 */ { rom[164], rom[165], rom[166], rom[167]} = 32'b100000_00000_00010_00000_00000000000;
  /* 33 */ { rom[168], rom[169], rom[170], rom[171]} = 32'b100000_00000_00011_00000_00000000001;
  /* 34 */ { rom[172], rom[173], rom[174], rom[175]} = 32'b100000_00000_01001_00000_00000000010;
  
            {rom[176], rom[177], rom[178], rom[179]} = 32'd0;
            {rom[180], rom[181], rom[182], rom[183]} = 32'd0;
            
  /* 35 */ {rom[184], rom[185], rom[186], rom[187]} = 32'b001010_00011_01001_01000_00000000000;
  
            {rom[188], rom[189], rom[190], rom[191]} = 32'd0; 
            {rom[192], rom[193], rom[194], rom[195]} = 32'd0; 
            
 /* 36 */   {rom[196], rom[197], rom[198], rom[199]} = 32'b000001_00100_01000_01000_00000000000;
 
            {rom[200], rom[201], rom[202], rom[203]} = 32'd0; 
            {rom[204], rom[205], rom[206], rom[207]} = 32'd0;
            
   /* 37 */ {rom[208], rom[209], rom[210], rom[211]} = 32'b100100_01000_00101_00000_00000000000;
           
            {rom[212], rom[213], rom[214], rom[215]} = 32'd0; 
            { rom[216], rom[217], rom[218], rom[219]} = 32'd0;

   /* 38 */ {rom[220], rom[221], rom[222], rom[223]} = 32'b100100_01000_00110_11111_11111111100; 
         
            {rom[224], rom[ 225], rom[226], rom[227]} = 32'd0; 
            {rom[228], rom[229], rom[230], rom[231]} = 32'd0;
            
   /* 39 */ {rom[232], rom[233], rom[234], rom[235]} = 32'b000011_00101_00110_01001_00000000000;
   /* 40 */ { rom[236], rom[237], rom[238], rom[239]} = 32'b100000_00000_01010_10000_00000000000;
   /* 41 */ { rom[240], rom[241], rom[242], rom[243]} = 32'b100000_00000_01011_00000_00000010000;
   
            {rom[244], rom[245], rom[246], rom[247]} = 32'd0; 
            {rom[248], rom[249], rom[250], rom[251]} = 32'd0;
            
   /* 42 */ {rom[252], rom[253], rom[254], rom[255]} = 32'b001010_01010_01011_01010_00000000000;
   
            {rom[256], rom[257], rom[258], rom[259]} = 32'd0; 
            { rom[260], rom[261], rom[262], rom[263]} = 32'd0;
            
   /* 43 */ { rom[264], rom[265], rom[266], rom[267]} = 32'b000101_01001_01010_01001_00000000000;
            { rom[268], rom[269], rom[270], rom[271]} = 32'd0; 
            { rom[272], rom[273], rom[274], rom[275]} = 32'd0;
   /* 44 */ { rom[276], rom[277], rom[278], rom[279]} = 32'b101000_01001_00000_00000_00000000010;
   /* 45 */ {rom[280], rom[281], rom[282], rom[283]} = 32'b100101_01000_00101_11111_11111111100;
   /* 46 */ {rom[284], rom[285], rom[286], rom[287]} = 32'b100101_01000_00110_00000_00000000000;
   /* 47 */ {rom[288], rom[289], rom[290], rom[291]} = 32'b100000_00011_00011_00000_00000000001;
   
             {rom[292], rom[293], rom[294], rom[295]} = 32'd0; 
             { rom[296], rom[297], rom[298], rom[299]} = 32'd0;
             
   /* 48 */ {rom[300], rom[301], rom[302], rom[303]}= 32'b101001_00001_00011_1111111111011110;
   /* 49 */ {rom[304], rom[305], rom[306], rom[307]} = 32'b100000_00010_00010_00000_00000000001;
   
            {rom[308], rom[309], rom[310], rom[311]} = 32'd0; 
            {rom[312], rom[313], rom[314], rom[315]} = 32'd0;
            
   /* 50 */ {rom[316], rom[317], rom[318], rom[319]} = 32'b101001_00001_00010_1111111111011001;
   /* 51 */ {rom[320], rom[321], rom[322], rom[323]} = 32'b100000_00000_00001_00000_10000000000;

            {rom[324], rom[325], rom[326], rom[327]} = 32'd0; 
            {rom[328], rom[329], rom[330], rom[331]} = 32'd0;
            
  /* 52 */ { rom[332], rom[333], rom[334], rom[335]} = 32'b100100_00001_00010_00000_00000000000;
   /* 53 */ { rom[336], rom[337], rom[338], rom[339]} = 32'b100100_00001_00011_00000_00000000100;
   /* 54 */{ rom[340], rom[341], rom[342], rom[343]} = 32'b100100_00001_00100_00000_00000001000;
   /* 55 */ { rom[344], rom[345], rom[346], rom[347]}= 32'b100100_00001_00100_00000_01000001000;
   /* 56 */{ rom[348], rom[349], rom[350], rom[351]} = 32'b100100_00001_00100_00000_10000001000;


/* 57 */ { rom[352], rom[353], rom[354], rom[355]}= 32'b100100_00001_00101_00000_00000001100;
/* 58 */  { rom[356], rom[357], rom[358], rom[359]}= 32'b100100_00001_00110_00000_00000010000;
/* 59 */ { rom[360], rom[361], rom[362], rom[363]}= 32'b100100_00001_00111_00000_00000010100;
/* 60 */  { rom[364], rom[365], rom[366], rom[367]}= 32'b100100_00001_01000_00000_00000011000;
/* 61 */ { rom[368], rom[369], rom[370], rom[371]} = 32'b100100_00001_01001_00000_00000011100;
/* 62 */ { rom[372], rom[373], rom[374], rom[375]}  = 32'b100100_00001_01010_00000_00000100000;
/* 63 */ { rom[376], rom[377], rom[378], rom[379]}= 32'b100100_00001_01011_00000_00000100100;
/* 64 */ { rom[380], rom[381], rom[382], rom[383]} = 32'b101010_00000_00000_11111_11111111111;


	 	end
  end
  
  assign instruction = (reset)? 32'd0 : {rom[address], rom[address+1], rom[address+2], rom[address+3]};

endmodule 